module ROB(clk, reset_n, );
    input clk, reset_n;
endmodule

module ROB_one(clk, reset_n, );