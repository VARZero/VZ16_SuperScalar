/*  ====================================
    VZ16(MMC16) Instruction Set Decoder
    ==================================== */

module scRenamer();
    input clk, reset_n;
    input [15:0] i0, i1, i2, i3;
    output 
endmodule
